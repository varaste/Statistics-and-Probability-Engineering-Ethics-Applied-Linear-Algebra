library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--
entity ROM is
	port(-- Address
				"0011",		-- 00
				"1100",		-- 01
				"0010",		-- 02
				"1000",		-- 03
				"1010",		-- 04
				
				"0010",		-- 27
				"0100",		-- 28
				"0110",		-- 29
				"1000",		-- 30
				"1010"		-- 

