ibrary IEEE;
use IEC;
        clk: in STD_LOGIC;
        clr: 
