entity logical_alu is
port ( a,b : in  std_logic_vector(3 downto 0);
       op : in  std_l
