

architecture dataflow of ha is
begin
    s<= a xor b ;
    co<= a and b ;
end;
