library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--
entity ROM is
	port(-- Address
				"0011",		-- 00
				"1100",		-- 01
				"0010",		-- 02
				"1000",		-- 03
				"1010",		-- 04
				"0010",		-- 05
				"1101",		-- 06
				"1100",		-- 07
				"1101",		-- 08
				"1110",		-- 09
				"0010",		-- 10
				"0100",		-- 11
			"1100",		-- 24
				"1110",		-- 25
				"0000",		-- 26
				"0010",		-- 27
				"0100",		-- 28
				"0110",		-- 29
				"1000",		-- 30
				"1010"		-- 

