library ieee;
use ieee.std_lclk)
     nt AND clk=
