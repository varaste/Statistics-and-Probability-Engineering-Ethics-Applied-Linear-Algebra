_arch of flipwait is
begink='1';
         q<=d;
   end process;      
end flipwait_arch;
