library IEEE;
use IEEE.std_logic_1164.all;

entity flipt is
    port (
        t,clk
arch
		else
		q<=q;
		end if;
	end if;
end process;
end flipt_arch;
