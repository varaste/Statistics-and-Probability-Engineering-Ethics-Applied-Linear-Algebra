
begin
	q <= signed(a) + signed(b);  	--(2)
end;
