ibrary IEEE;
use IEC;
