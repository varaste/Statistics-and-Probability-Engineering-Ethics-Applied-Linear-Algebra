library IEEE;
use IEEE.std_logic_1164.all;

entity registd is
        q: out STD_LOG
end registd_arch;
