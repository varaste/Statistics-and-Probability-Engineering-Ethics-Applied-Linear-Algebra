--
--*******Defining  and using function******

library ieee;
use ieee.std_logic_1164.all;
entity fu std
