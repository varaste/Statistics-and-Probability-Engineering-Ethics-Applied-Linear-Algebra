--
--*******Defining  and using function******
