library ieee;
use ieee.std_l
    begin
counter:process(clk)
     nt AND clk='1')then
		 cnt:=cnt+1;				--(2)
		 end if;
		count<=cnt;
		end process;
end;
