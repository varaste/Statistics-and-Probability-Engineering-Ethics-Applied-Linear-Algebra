library ieee;
use ieee.std_l
    begin
counter:process(clk)
     nt AND clk=
