--
--multiplexer 4 to 1 (4 bits), using 'with-- select' 
--
library IEEE;

architecture maxwith_arch of maxwith is
begin
