

    s<= a xor b ;
    co<= a and b ;
end;
