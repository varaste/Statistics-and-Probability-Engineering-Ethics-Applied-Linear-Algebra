library IEEE
          begin
            if reset='1' then
               cnt<=(others=>'0');
               elsif set='1' then
              end if;
end process count ;      
end counter1_arch;
